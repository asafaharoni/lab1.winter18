X_start_inst : X_start PORT MAP (
		result	 => result_sig
	);
